`timescale 1ns / 1ps

module alu_tb;
  integer SIZE 7;

  reg[SIZE:0] a, b;
  reg[1:0] sel;

  
endmodule
